// ----  Probes  ----
`define PROBE_F_PC      probe_f_pc
`define PROBE_F_INSN    probe_f_insn

`define PROBE_D_PC      probe_d_pc
`define PROBE_D_OPCODE  probe_d_opcode_o
`define PROBE_D_RD      probe_d_rd_o
`define PROBE_D_FUNCT3  probe_d_funct3
`define PROBE_D_RS1     probe_d_rs1_o
`define PROBE_D_RS2     probe_d_rs2_o
`define PROBE_D_FUNCT7  probe_d_funct7
`define PROBE_D_IMM     probe_d_imm_o
`define PROBE_D_SHAMT   probe_d_shamt_o
// ----  Probes  ----

// ----  Top module  ----
`define TOP_MODULE  pd2
// ----  Top module  ----

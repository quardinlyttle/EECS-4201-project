// ----  Probes  ----
`define PROBE_ADDR          probe_addr
`define PROBE_DATA_IN       probe_data_in
`define PROBE_DATA_OUT      probe_data_out
`define PROBE_READ_EN       probe_read_en
`define PROBE_WRITE_EN      probe_write_en

`define PROBE_F_PC          probe_f_pc
`define PROBE_F_INSN        probe_f_insn
// ----  Probes  ----

// ----  Top module  ----
`define TOP_MODULE          pd1
// ----  Top module  ----

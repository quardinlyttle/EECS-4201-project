// ----  Probes  ----
`define PROBE_ASSIGN_XOR_OP1 assign_xor_op1
`define PROBE_ASSIGN_XOR_OP2 assign_xor_op2
`define PROBE_ASSIGN_XOR_RES assign_xor_res

// Define other probes as required....
`define PROBE_ALU_OP1 assign_ALU_op1
`define PROBE_ALU_OP2 assign_ALU_op2
`define PROBE_ALU_RES assign_ALU_res
`define PROBE_ALU_SEL assign_ALU_sel
`define PROBE_ALU_NFLAG assign_ALU_nflag
`define PROBE_ALU_ZFLAG assign_ALU_zflag

`define PROBE_REG_IN  assign_reg_in
`define PROBE_REG_OUT assign_reg_out

`define PROBE_TSP_OP1 assign_TSP_op1
`define PROBE_TSP_OP2 assign_TSP_op2
`define PROBE_TSP_RES assign_TSP_res
// ----  Probes  ----

// ----  Top module  ----
`define TOP_MODULE  pd0
// ----  Top module  ----
